// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// File Name: cl_irq_up.v

`timescale 100ps/10ps 
`include "simulate_x_tick.vh"
`timescale 100ps/10ps 
`include "simulate_x_tick.vh"
module cl_irq_up (
   clk        //|< i
  ,irq        //|< i
  ,irq_ack    //|< i
  ,irq_pop    //|< i
  ,reset_     //|< i
  ,irq_req    //|> o
  ,irq_status //|> o
  );

input         clk;
input  [15:0] irq;
input  [15:0] irq_ack;
input  [15:0] irq_pop;
input         reset_;
output [15:0] irq_req;
output [15:0] irq_status;
wire   [15:0] irq_sync;



//// generated by ::sync -type 3D -inst irq_sync -input irq -output irq_sync -clock clk -reset reset_ -width 16

wire   [15:0] sync_ibus_0;
wire   [15:0] sync_rbus_0;
wire   [15:0] sync_bbus_0;
wire   [15:0] sync_sbus_0;

`undef SYNC_PL_NOSYNTHESIS_NOSYNTH_GCS
`ifndef SYNC_PL_NO_RANDOMIZATION
`ifndef SYNTH_LEVEL1_COMPILE
`ifndef SYNTHESIS
    `define SYNC_PL_NOSYNTHESIS_NOSYNTH_GCS
`endif
`endif
`endif

// VCS coverage off

`ifdef  SYNC_PL_NOSYNTHESIS_NOSYNTH_GCS
reg [15:0] RandSyncBusPipe_0 [0:1];
reg [15:0] RandSyncBusCurr_0;
reg [15:0] RandSyncBusNext_0;
reg [15:0] RandSyncBusRand_0;
reg [15:0] RandSyncBusPick_0;
reg [1:1] RandSyncBusKnown_0;
reg [1:1] RandSyncBusDelta_0;
reg        RandSyncEnable_0;
reg        RandSyncBusEnable_0;
reg        RandSyncBitEnable_0;
reg        RandSyncDiff_0;
reg        RandSyncDone_0;
reg        RandSyncSnap_0;
`endif
// VCS coverage on

// input bus

assign sync_ibus_0 = irq[15:0];

// random bus

`ifdef SYNC_PL_NOSYNTHESIS_NOSYNTH_GCS
  assign sync_rbus_0 = RandSyncBusRand_0;
`else 
  assign sync_rbus_0 = sync_ibus_0;
`endif

// buffer bus

assign sync_bbus_0 = sync_rbus_0;

 // sync bus


sync3d_c_ppp irq_sync_0 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[0]),
  .q(sync_sbus_0[0])
  );

sync3d_c_ppp irq_sync_1 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[1]),
  .q(sync_sbus_0[1])
  );

sync3d_c_ppp irq_sync_2 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[2]),
  .q(sync_sbus_0[2])
  );

sync3d_c_ppp irq_sync_3 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[3]),
  .q(sync_sbus_0[3])
  );

sync3d_c_ppp irq_sync_4 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[4]),
  .q(sync_sbus_0[4])
  );

sync3d_c_ppp irq_sync_5 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[5]),
  .q(sync_sbus_0[5])
  );

sync3d_c_ppp irq_sync_6 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[6]),
  .q(sync_sbus_0[6])
  );

sync3d_c_ppp irq_sync_7 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[7]),
  .q(sync_sbus_0[7])
  );

sync3d_c_ppp irq_sync_8 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[8]),
  .q(sync_sbus_0[8])
  );

sync3d_c_ppp irq_sync_9 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[9]),
  .q(sync_sbus_0[9])
  );

sync3d_c_ppp irq_sync_10 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[10]),
  .q(sync_sbus_0[10])
  );

sync3d_c_ppp irq_sync_11 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[11]),
  .q(sync_sbus_0[11])
  );

sync3d_c_ppp irq_sync_12 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[12]),
  .q(sync_sbus_0[12])
  );

sync3d_c_ppp irq_sync_13 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[13]),
  .q(sync_sbus_0[13])
  );

sync3d_c_ppp irq_sync_14 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[14]),
  .q(sync_sbus_0[14])
  );

sync3d_c_ppp irq_sync_15 (
  .clk(clk), 
  .clr_(reset_),
  .d(sync_bbus_0[15]),
  .q(sync_sbus_0[15])
  );

// defeating sync randomizer
`ifndef NO_PLI_OR_EMU
`ifndef GATES
`ifdef SYNC_PL_NOSYNTHESIS_NOSYNTH_GCS

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_0.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_0.first_stage_of_sync.mode = 0;
`endif

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_1.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_1.first_stage_of_sync.mode = 0;
`endif

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_2.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_2.first_stage_of_sync.mode = 0;
`endif

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_3.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_3.first_stage_of_sync.mode = 0;
`endif

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_4.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_4.first_stage_of_sync.mode = 0;
`endif

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_5.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_5.first_stage_of_sync.mode = 0;
`endif

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_6.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_6.first_stage_of_sync.mode = 0;
`endif

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_7.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_7.first_stage_of_sync.mode = 0;
`endif

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_8.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_8.first_stage_of_sync.mode = 0;
`endif

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_9.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_9.first_stage_of_sync.mode = 0;
`endif

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_10.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_10.first_stage_of_sync.mode = 0;
`endif

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_11.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_11.first_stage_of_sync.mode = 0;
`endif

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_12.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_12.first_stage_of_sync.mode = 0;
`endif

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_13.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_13.first_stage_of_sync.mode = 0;
`endif

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_14.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_14.first_stage_of_sync.mode = 0;
`endif

`ifdef NVTOOLS_SYNC2D_GENERIC_CELL
  defparam irq_sync_15.NV_GENERIC_CELL.first_stage_of_sync.mode = 0;
`else
  defparam irq_sync_15.first_stage_of_sync.mode = 0;
`endif

`endif
`endif
`endif

// output bus

assign irq_sync = sync_sbus_0;

// VCS coverage off
`ifndef NO_PLI_OR_EMU
`ifdef SYNC_PL_NOSYNTHESIS_NOSYNTH_GCS

initial begin
  if ($test$plusargs("RandSyncInfo")) $display ("INFO: RandSync:  @ %m");
end

initial begin
  RandSyncEnable_0 = 1'b1;
  if ($test$plusargs("RandSyncGlobalDisable")) RandSyncEnable_0 = 1'b0;
  if ($test$plusargs("RandSyncLocalDisable")) RandSyncEnable_0 = 1'b0;
end

// SRC before DSTCLK: new SRC is sampled to CUR, CUR is sampled to PRE, CUR/PRE are randomized.
// SRC equals DSTCLK: new SRC is sampled to CUR, CUR is sampled to PRE, CUR/PRE are randomized.
// SRC after  DSTCLK: old SRC is sampled again to CUR (NOP), CUR is sampled to PRE, CUR == PRE.

// curr (glitch filter)
always @(sync_ibus_0) begin
  RandSyncBusCurr_0 <= sync_ibus_0;
end

// snap
initial RandSyncSnap_0 = 1'b0;
always @(posedge clk) begin 
  RandSyncSnap_0 <= (RandSyncSnap_0 === 1'bx)? 1'b0 : !RandSyncSnap_0; 
end

// eval
always @(RandSyncBusCurr_0 or RandSyncSnap_0 or negedge reset_) begin : rand_sync_block_0
  integer i, j;

  // bump
  for (i=1; i>=1; i=i-1) begin
    RandSyncBusPipe_0[i] = RandSyncBusPipe_0[i-1];
  end
  RandSyncBusPipe_0[0] = RandSyncBusCurr_0; 
 
  // next
  RandSyncBusNext_0 = RandSyncBusPipe_0[0]; 
 
  // rand 
  if (RandSyncEnable_0 && reset_) begin
    // known
    for (i=1; i>=1; i=i-1) begin
      RandSyncBusKnown_0[i] = |RandSyncBusPipe_0[i] !== 1'bx;
    end
    // delta
    for (i=1; i>=1; i=i-1) begin
      RandSyncBusDelta_0[i] = |(RandSyncBusPipe_0[i] ^ RandSyncBusPipe_0[i-1]);
    end
    if (&RandSyncBusKnown_0 && |RandSyncBusDelta_0) begin 
      RandSyncBusNext_0 = RandSyncBusPipe_0[1]; 
      RandSyncBusEnable_0 = prand_inst0(1, 100) > (100 - 50);
      if (RandSyncBusEnable_0) begin 
        RandSyncDone_0 = 1'b0;
        for (i=1; i>=1; i=i-1) begin
          RandSyncDiff_0 = RandSyncBusPipe_0[i] !== RandSyncBusPipe_0[i-1];
          if (RandSyncDiff_0 && !RandSyncDone_0) begin
            RandSyncBusPickTask_0 (RandSyncBusPipe_0[i], RandSyncBusPipe_0[i-1]);
            if (RandSyncBusNext_0 !== RandSyncBusPick_0) begin
              RandSyncBusNext_0 = RandSyncBusPick_0;
              RandSyncDone_0 = 1'b1;
            end
          end
        end
      end
    end
  end
  RandSyncBusRand_0 = RandSyncBusNext_0;
end

// task
task RandSyncBusPickTask_0; // rand value = mixture
  input [15:0] RandSyncTaskBusPrev_0;
  input [15:0] RandSyncTaskBusCurr_0;
  integer i;
  for (i=0; i<=15; i=i+1) begin
    if (RandSyncTaskBusCurr_0[i] === RandSyncTaskBusPrev_0[i]) begin
      RandSyncBusPick_0[i] = RandSyncTaskBusCurr_0[i];
    end else begin
      RandSyncBitEnable_0 = prand_inst1(1, 100) > (100 - 50);
      RandSyncBusPick_0[i] = (RandSyncBitEnable_0)? RandSyncTaskBusCurr_0[i] : RandSyncTaskBusPrev_0[i];
    end
  end
endtask


`ifdef SYNTH_LEVEL1_COMPILE
`else
`ifdef SYNTHESIS
`else
`ifdef PRAND_VERILOG
// Only verilog needs any local variables
reg [47:0] prand_local_seed0;
reg prand_initialized0;
reg prand_no_rollpli0;
`endif
`endif
`endif

function [31:0] prand_inst0;
//VCS coverage off
    input [31:0] min;
    input [31:0] max;
    reg [32:0] diff;
    
    begin
`ifdef SYNTH_LEVEL1_COMPILE
        prand_inst0 = min;
`else
`ifdef SYNTHESIS
        prand_inst0 = min;
`else
`ifdef PRAND_VERILOG
        if (prand_initialized0 !== 1'b1) begin
            prand_no_rollpli0 = $test$plusargs("NO_ROLLPLI");
            if (!prand_no_rollpli0)
                prand_local_seed0 = {$prand_get_seed(0), 16'b0};
            prand_initialized0 = 1'b1;
        end
        if (prand_no_rollpli0) begin
            prand_inst0 = min;
        end else begin
            diff = max - min + 1;
            prand_inst0 = min + prand_local_seed0[47:16] % diff;
            // magic numbers taken from Java's random class (same as lrand48)
            prand_local_seed0 = prand_local_seed0 * 48'h5deece66d + 48'd11;
        end
`else
`ifdef PRAND_OFF
        prand_inst0 = min;
`else
        prand_inst0 = $RollPLI(min, max, "auto");
`endif
`endif
`endif
`endif
    end
//VCS coverage on
endfunction


`ifdef SYNTH_LEVEL1_COMPILE
`else
`ifdef SYNTHESIS
`else
`ifdef PRAND_VERILOG
// Only verilog needs any local variables
reg [47:0] prand_local_seed1;
reg prand_initialized1;
reg prand_no_rollpli1;
`endif
`endif
`endif

function [31:0] prand_inst1;
//VCS coverage off
    input [31:0] min;
    input [31:0] max;
    reg [32:0] diff;
    
    begin
`ifdef SYNTH_LEVEL1_COMPILE
        prand_inst1 = min;
`else
`ifdef SYNTHESIS
        prand_inst1 = min;
`else
`ifdef PRAND_VERILOG
        if (prand_initialized1 !== 1'b1) begin
            prand_no_rollpli1 = $test$plusargs("NO_ROLLPLI");
            if (!prand_no_rollpli1)
                prand_local_seed1 = {$prand_get_seed(1), 16'b0};
            prand_initialized1 = 1'b1;
        end
        if (prand_no_rollpli1) begin
            prand_inst1 = min;
        end else begin
            diff = max - min + 1;
            prand_inst1 = min + prand_local_seed1[47:16] % diff;
            // magic numbers taken from Java's random class (same as lrand48)
            prand_local_seed1 = prand_local_seed1 * 48'h5deece66d + 48'd11;
        end
`else
`ifdef PRAND_OFF
        prand_inst1 = min;
`else
        prand_inst1 = $RollPLI(min, max, "auto");
`endif
`endif
`endif
`endif
    end
//VCS coverage on
endfunction


`endif
`endif
// VCS coverage on


cl_irq_up_bit CL_IRQ_UP_BIT0 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[0])      //|< i
  ,.irq_in     (irq_sync[0])     //|< w
  ,.irq_pop    (irq_pop[0])      //|< i
  ,.irq_req    (irq_req[0])      //|> o
  ,.irq_status (irq_status[0])   //|> o
  );

cl_irq_up_bit CL_IRQ_UP_BIT1 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[1])      //|< i
  ,.irq_in     (irq_sync[1])     //|< w
  ,.irq_pop    (irq_pop[1])      //|< i
  ,.irq_req    (irq_req[1])      //|> o
  ,.irq_status (irq_status[1])   //|> o
  );

cl_irq_up_bit CL_IRQ_UP_BIT2 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[2])      //|< i
  ,.irq_in     (irq_sync[2])     //|< w
  ,.irq_pop    (irq_pop[2])      //|< i
  ,.irq_req    (irq_req[2])      //|> o
  ,.irq_status (irq_status[2])   //|> o
  );

cl_irq_up_bit CL_IRQ_UP_BIT3 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[3])      //|< i
  ,.irq_in     (irq_sync[3])     //|< w
  ,.irq_pop    (irq_pop[3])      //|< i
  ,.irq_req    (irq_req[3])      //|> o
  ,.irq_status (irq_status[3])   //|> o
  );

cl_irq_up_bit CL_IRQ_UP_BIT4 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[4])      //|< i
  ,.irq_in     (irq_sync[4])     //|< w
  ,.irq_pop    (irq_pop[4])      //|< i
  ,.irq_req    (irq_req[4])      //|> o
  ,.irq_status (irq_status[4])   //|> o
  );

cl_irq_up_bit CL_IRQ_UP_BIT5 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[5])      //|< i
  ,.irq_in     (irq_sync[5])     //|< w
  ,.irq_pop    (irq_pop[5])      //|< i
  ,.irq_req    (irq_req[5])      //|> o
  ,.irq_status (irq_status[5])   //|> o
  );

cl_irq_up_bit CL_IRQ_UP_BIT6 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[6])      //|< i
  ,.irq_in     (irq_sync[6])     //|< w
  ,.irq_pop    (irq_pop[6])      //|< i
  ,.irq_req    (irq_req[6])      //|> o
  ,.irq_status (irq_status[6])   //|> o
  );

cl_irq_up_bit CL_IRQ_UP_BIT7 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[7])      //|< i
  ,.irq_in     (irq_sync[7])     //|< w
  ,.irq_pop    (irq_pop[7])      //|< i
  ,.irq_req    (irq_req[7])      //|> o
  ,.irq_status (irq_status[7])   //|> o
  );

cl_irq_up_bit CL_IRQ_UP_BIT8 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[8])      //|< i
  ,.irq_in     (irq_sync[8])     //|< w
  ,.irq_pop    (irq_pop[8])      //|< i
  ,.irq_req    (irq_req[8])      //|> o
  ,.irq_status (irq_status[8])   //|> o
  );

cl_irq_up_bit CL_IRQ_UP_BIT9 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[9])      //|< i
  ,.irq_in     (irq_sync[9])     //|< w
  ,.irq_pop    (irq_pop[9])      //|< i
  ,.irq_req    (irq_req[9])      //|> o
  ,.irq_status (irq_status[9])   //|> o
  );

cl_irq_up_bit CL_IRQ_UP_BIT10 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[10])     //|< i
  ,.irq_in     (irq_sync[10])    //|< w
  ,.irq_pop    (irq_pop[10])     //|< i
  ,.irq_req    (irq_req[10])     //|> o
  ,.irq_status (irq_status[10])  //|> o
  );

cl_irq_up_bit CL_IRQ_UP_BIT11 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[11])     //|< i
  ,.irq_in     (irq_sync[11])    //|< w
  ,.irq_pop    (irq_pop[11])     //|< i
  ,.irq_req    (irq_req[11])     //|> o
  ,.irq_status (irq_status[11])  //|> o
  );

cl_irq_up_bit CL_IRQ_UP_BIT12 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[12])     //|< i
  ,.irq_in     (irq_sync[12])    //|< w
  ,.irq_pop    (irq_pop[12])     //|< i
  ,.irq_req    (irq_req[12])     //|> o
  ,.irq_status (irq_status[12])  //|> o
  );

cl_irq_up_bit CL_IRQ_UP_BIT13 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[13])     //|< i
  ,.irq_in     (irq_sync[13])    //|< w
  ,.irq_pop    (irq_pop[13])     //|< i
  ,.irq_req    (irq_req[13])     //|> o
  ,.irq_status (irq_status[13])  //|> o
  );

cl_irq_up_bit CL_IRQ_UP_BIT14 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[14])     //|< i
  ,.irq_in     (irq_sync[14])    //|< w
  ,.irq_pop    (irq_pop[14])     //|< i
  ,.irq_req    (irq_req[14])     //|> o
  ,.irq_status (irq_status[14])  //|> o
  );

cl_irq_up_bit CL_IRQ_UP_BIT15 (
   .clk        (clk)             //|< i
  ,.reset_     (reset_)          //|< i
  ,.irq_ack    (irq_ack[15])     //|< i
  ,.irq_in     (irq_sync[15])    //|< w
  ,.irq_pop    (irq_pop[15])     //|< i
  ,.irq_req    (irq_req[15])     //|> o
  ,.irq_status (irq_status[15])  //|> o
  );


endmodule // cl_irq_up


